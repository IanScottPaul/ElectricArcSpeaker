module EAS(input logic clk, rx, RTS, output logic tx, CTS, )